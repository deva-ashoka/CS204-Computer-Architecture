// Not Circuit - Assignment 1 - Q1 Figure 0 - A_bar

module andCircuit (A, A_bar);

input A;
output A_bar;

not not1(A_bar, A);

endmodule
