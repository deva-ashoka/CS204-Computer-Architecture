// Or Circuit - Assignment 1 - Q1 Figure 0 - A or B

module andCircuit (A, B, AorB);

input A, B;
output AorB;

or or1(AorB, A, B);

endmodule
