//inverter logic gate - created by Deva

module inverter (
input1,
output1
);

input input1;
output output1;

assign output1 = ~ input1;

endmodule
