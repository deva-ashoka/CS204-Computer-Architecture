// And Circuit - Assignment 1 - Q1 Figure 0 - AB

module andCircuit (A, B, AB);

input A, B;
output AB;

and and1(AB, A, B);

endmodule
